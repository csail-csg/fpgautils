
// Copyright (c) 2017 Massachusetts Institute of Technology
// 
// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.
// 
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

import ResetGuard::*;

// some xilinx IP automatically reset
// we wait several cycles to make sure the reset completes
// we also block signals on the IP before reset of current clock domain completes
// because such signals may be garbage

interface WaitAutoReset#(numeric type logCycles);
    method Bool isReady;
endinterface

module mkWaitAutoReset(WaitAutoReset#(logCycles));
    Reg#(Bit#(logCycles)) cnt <- mkReg(0);
    Reg#(Bool) init <- mkReg(False);
    
    ResetGaurd rg <- mkResetGuard;

    rule doInit(!init);
        cnt <= cnt + 1;
        if(cnt == maxBound) begin
            init <= True;
        end
    endrule

    method Bool isReady;
        return init && rg.isReady;
    endmethod
endmodule
